
module pong
	(
		CLOCK_50,						//	On Board 50 MHz
	);
